
////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:    16:31:33 09/14/09
// Design Name:    
// Module Name:    and_gate_2input
// Project Name:   
// Target Device:  
// Tool versions:  
// Description:
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////
module and_gate_2input(a, b, y);
    input a;
    input b;
    output y;

	 assign y = a & b ;

endmodule